library verilog;
use verilog.vl_types.all;
entity mach_test is
end mach_test;
