library verilog;
use verilog.vl_types.all;
entity M2_test is
end M2_test;
