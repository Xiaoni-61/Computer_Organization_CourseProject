library verilog;
use verilog.vl_types.all;
entity DM_test is
end DM_test;
