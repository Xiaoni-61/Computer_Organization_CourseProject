library verilog;
use verilog.vl_types.all;
entity im_test is
end im_test;
