library verilog;
use verilog.vl_types.all;
entity EXT_test is
end EXT_test;
