library verilog;
use verilog.vl_types.all;
entity mips_test is
end mips_test;
