library verilog;
use verilog.vl_types.all;
entity GPR_test is
end GPR_test;
