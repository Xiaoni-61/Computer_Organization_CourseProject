library verilog;
use verilog.vl_types.all;
entity ifu_test is
end ifu_test;
