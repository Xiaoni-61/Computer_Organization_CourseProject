module ALUtoDM_addr(ALUout,addr);
  input [31:0] ALUout;
  output [9:0] addr;
  
  assign addr={ALUout[9:0]};
  
endmodule
