library verilog;
use verilog.vl_types.all;
entity ALU_test is
end ALU_test;
