module ifu(clk,reset,jsome,jr,npc_sel,zero,pcc,AOut,code,enpc);      //pcc is for jal, AOut is for jr
  input enpc;
  input clk,reset,npc_sel,zero;
  
  input jsome;
  input jr;
  input [31:0] AOut;
  output [31:0] code;
  
  output reg [31:0]pcc;
  
  wire [31:0] t1,t0,extout,temp;              //wire?????
  reg [31:0] pcnew,pc;
  wire [15:0] imm;
  
  
  
  im_1k im1(.addr(pc[9:0]),.dout(code));
  
  //assign insout={im[pc[9:0]],im[pc[9:0]+1],im[pc[9:0]+2],im[pc[9:0]+3]};    //for getting imm16
  assign imm=code[15:0];
  assign temp={{16{imm[15]}},imm};
  assign extout=temp<<2;
  //assign pcc=pc+4;
  
  always@(posedge clk)
  begin
    if(jsome)
      pcnew={pc[31:28],code[25:0],{2{1'b0}}};
    else if(npc_sel&&zero)
      pcnew=t1;
    else if(jr)
      pcnew=AOut;
    
    else
      pcnew=t0;
      
      pcc=pc+4;
  end
  
  always@(posedge clk,posedge reset)
  begin
    if(reset) pc=32'h0000_3000;
    else
      if(enpc)
      pc=pcnew;
  end
  
  
  assign t0=pc+4;
  assign t1=t0+extout;
 
endmodule
