library verilog;
use verilog.vl_types.all;
entity M1_test is
end M1_test;
